
*The Complete pixel sensor
.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS


XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

XC1 VCMP_OUT VSTORE VRAMP VDD VSS COMP

XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS

*Memory bank, ready made
.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS

*Memory cell, ready made
.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS

*Actual photogate, ready i think
.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

* Capacitor to model gate-source capacitance
C1 VSTORE VSS 100f
Rleak VSTORE VSS 100T

* Switch to reset voltage on capacitor
BR1 VRESET VSTORE I=V(ERASE)*V(VRESET,VSTORE)/1k

* Switch to expose pixel
BR2 VPG VSTORE I=V(EXPOSE)*V(VSTORE,VPG)/1k

* Model photocurrent
Rphoto VPG VSS 1G
.ENDS

*Comparator
.SUBCKT COMP VCMP_OUT VSTORE VRAMP VDD VSS

*Can be tuned
VBIAS1 VBIAS1 VSS dc 0.9
VBIAS2 VBIAS2 VSS dc 0.65

*Transistor widths can be tuned

*Diff pair
M1 VG1 VG1 VDD VDD pmos w=1u l=0.13u
M2 VCMP VG1 VDD VDD pmos w=1u l=0.13u
M3 VG1 VSTORE VC VC nmos w=0.5u l=0.13u
M4 VCMP VRAMP VC VC nmos w=0.5u l=0.13u
M7 VCMP_INV VCMP VDD VDD pmos w=1.2u l=0.13u

*Current mirror
M5 VC VBIAS1 VSS VSS nmos w=0.5u l=0.13u
M6 VCMP_INV VBIAS2 VSS VSS nmos w=0.5u l=0.13u

*Inverter
M8 VCMP_OUT VCMP_INV VDD VDD pmos w=1.2u l=0.13u
M9 VCMP_OUT VCMP_INV VSS VSS nmos W=0.5u l=0.13u

.ENDS
